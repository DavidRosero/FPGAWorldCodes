library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.std_logic_arith.all;
USE WORK.COMANDOS_LCD_REVC.ALL;

entity LIB_LCD_INTESC_REVC is


PORT(CLK: IN STD_LOGIC;

-------------------------------------------------------
-------------PUERTOS DE LA LCD (NO BORRAR)-------------
	  RS : OUT STD_LOGIC;									  --
	  RW : OUT STD_LOGIC;									  --
	  ENA : OUT STD_LOGIC;									  --
	  CORD : IN STD_LOGIC;									  --
	  CORI : IN STD_LOGIC;									  --
	  DATA_LCD: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);     --
	  BLCD :  OUT STD_LOGIC_VECTOR(7 DOWNTO 0);       --
-------------------------------------------------------
	  
-----------------------------------------------------------
--------------ABAJO ESCRIBE TUS PUERTOS--------------------	
		ECO : IN STD_LOGIC;
		TRIGGER : OUT STD_LOGIC;
		DATO_LISTO : OUT STD_LOGIC
	  );



end LIB_LCD_INTESC_REVC;

architecture Behavioral of LIB_LCD_INTESC_REVC is

-----------------------------------------------------------------
---------------SE�ALES DE LA LCD (NO BORRAR)---------------------
TYPE RAM IS ARRAY (0 TO  60) OF STD_LOGIC_VECTOR(8 DOWNTO 0);  --
																					--
SIGNAL INST : RAM;													--
																					--
COMPONENT PROCESADOR_LCD_REVC is											--
																					--
PORT(CLK : IN STD_LOGIC;													--
	  VECTOR_MEM : IN STD_LOGIC_VECTOR(8 DOWNTO 0);					--
	  INC_DIR : OUT INTEGER RANGE 0 TO 1024;							--
	  CORD : IN STD_LOGIC;													--
	  CORI : IN STD_LOGIC;													--
	  RS : OUT STD_LOGIC;													--
	  RW : OUT STD_LOGIC;													--
	  DELAY_COR : IN INTEGER RANGE 0 TO 1000;							--
	  BD_LCD : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);			         --
	  ENA  : OUT STD_LOGIC;													--
	  C1A,C2A,C3A,C4A : IN STD_LOGIC_VECTOR(39 DOWNTO 0);       --
	  C5A,C6A,C7A,C8A : IN STD_LOGIC_VECTOR(39 DOWNTO 0);       --
	  DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)							--
		);																			--
																					--
end  COMPONENT PROCESADOR_LCD_REVC;	
-------------------------
COMPONENT INTESC_LIB_ULTRASONICO_RevC is

PORT(
		CLK 			 : IN  STD_LOGIC;                   -- Reloj del FPGA.
		ECO 			 : IN  STD_LOGIC;                   -- Eco del sensor ultras�nico.
		TRIGGER 		 : OUT STD_LOGIC;                   -- Trigger del sensor ultras�nico.
		DATO_LISTO 	 : OUT STD_LOGIC;                   -- Bandera que indica cuando el valor de la distancia es correcto.
		DISTANCIA_CM : OUT STD_LOGIC_VECTOR(8 DOWNTO 0) -- Valor de la distancia en cent�metros-
);

end COMPONENT INTESC_LIB_ULTRASONICO_RevC;
------------------------
									--
																					--
COMPONENT CARACTERES_ESPECIALES_REVC is										--
																					--
PORT( C1,C2,C3,C4:OUT STD_LOGIC_VECTOR(39 DOWNTO 0);				--
		C5,C6,C7,C8:OUT STD_LOGIC_VECTOR(39 DOWNTO 0);				--
		CLK : IN STD_LOGIC													--
		);																			--
																					--
end COMPONENT CARACTERES_ESPECIALES_REVC;	

             								--


                  							--

																					--
CONSTANT CHAR1 : INTEGER := 1;											--
CONSTANT CHAR2 : INTEGER := 2;											--
CONSTANT CHAR3 : INTEGER := 3;											--
CONSTANT CHAR4 : INTEGER := 4;											--
CONSTANT CHAR5 : INTEGER := 5;											--
CONSTANT CHAR6 : INTEGER := 6;											--
CONSTANT CHAR7 : INTEGER := 7;											--
CONSTANT CHAR8 : INTEGER := 8;											--
																					--
																					--
SIGNAL DIR : INTEGER RANGE 0 TO 1024 := 0;							--
SIGNAL VECTOR_MEM_S : STD_LOGIC_VECTOR(8 DOWNTO 0);				--
SIGNAL RS_S, RW_S, E_S : STD_LOGIC;										--
SIGNAL DATA_S : STD_LOGIC_VECTOR(7 DOWNTO 0);						--
SIGNAL DIR_S : INTEGER RANGE 0 TO 1024;								--
SIGNAL DELAY_COR : INTEGER RANGE 0 TO 1000;							--
SIGNAL C1S,C2S,C3S,C4S : STD_LOGIC_VECTOR(39 DOWNTO 0);	      --
SIGNAL C5S,C6S,C7S,C8S : STD_LOGIC_VECTOR(39 DOWNTO 0);  	   --
----------------------------------------------------------------
-----------------------------------------------------------------


---------------------------------------------------------
--------------AGREGA TUS SE�ALES AQU�--------------------
SIGNAL DISTANCIA_CM : STD_LOGIC_VECTOR(8 DOWNTO 0);
--SIGNAL DISTANCIA_CM0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL DISTANCIA_CM1 : INTEGER RANGE 0 TO 999;
SIGNAL CENTENAS,DECENAS,UNIDADES :INTEGER RANGE 0 TO 9 :=0;
---------------------------------------------------------

BEGIN
--
process(DISTANCIA_CM)
  begin
    DISTANCIA_CM1 <= TO_INTEGER(UNSIGNED(DISTANCIA_CM));
  end process;



-----------------------------------------------------------
------------COMPONENTES PARA LCD (NO BORRAR)---------------
U1 : PROCESADOR_LCD_REVC PORT MAP(CLK  => CLK,				--
									 VECTOR_MEM => VECTOR_MEM_S,	--
									 RS  => RS_S,						--
									 RW  => RW_S,						--
									 ENA => E_S,						--
									 INC_DIR => DIR_S,				--
									 DELAY_COR => DELAY_COR,		--
									 BD_LCD => BLCD,					--
									 CORD => CORD,						--
									 CORI => CORI,						--
									 C1A =>C1S,  					   --	
									 C2A =>C2S,							--
									 C3A =>C3S,							--
									 C4A =>C4S,							--
									 C5A =>C5S,							--
									 C6A =>C6S,							--
									 C7A =>C7S,							--
									 C8A =>C8S,							--
									 DATA  => DATA_S );				--
																			--
U2 : CARACTERES_ESPECIALES_REVC PORT MAP(C1 =>C1S,			--	
									C2 =>C2S,							--
									C3 =>C3S,							--
									C4 =>C4S,							--
									C5 =>C5S,							--
									C6 =>C6S,							--
									C7 =>C7S,						   --
									C8 =>C8S,							--
									CLK => CLK							--
									);	
U3:INTESC_LIB_ULTRASONICO_RevC PORT MAP(CLK => CLK,
													 ECO => ECO,
													 TRIGGER => TRIGGER,
													 DATO_LISTO => DATO_LISTO,
													 DISTANCIA_CM => DISTANCIA_CM
														);									
																			--
DIR <= DIR_S;															--
VECTOR_MEM_S <= INST(DIR);								--
																			--
RS <= RS_S;																--
RW <= RW_S;																--
ENA <= E_S;																--
DATA_LCD <= DATA_S;

																			--
													                  --
-----------------------------------------------------------


DELAY_COR <= 600; --Modificar esta variable para la velocidad del corrimiento.

-------------------------------------------------------------------
-----------------ABAJO ESCRIBE TU C�DIGO EN VHDL-------------------

CENTENAS <= DISTANCIA_CM1 / 100;
DECENAS <= (DISTANCIA_CM1/10) MOD 10;
UNIDADES <= DISTANCIA_CM1 MOD 10;
-----------------------------------------------------------------------------------------
-------------------------ABAJO ESCRIBE TU C�DIGO PARA LA LCD-----------------------------

INST(0) <= LCD_INI("00");

INST(1) <= CHAR(MD);
INST(2) <= CHAR(I);
INST(3) <= CHAR(S);
INST(4) <= CHAR(T);
INST(5) <= CHAR(A);
INST(6) <= CHAR(N);
INST(7) <= CHAR(C);
INST(8) <= CHAR(I);
INST(9) <= CHAR(A);
INST(10) <= CHAR_ASCII(X"3A");

INST(11) <= BUCLE_INI(1);

INST(12) <= POS(2,2);
INST(13) <= INT_NUM(CENTENAS);

INST(14) <= POS(2,3);
INST(15) <= INT_NUM(DECENAS);

INST(16) <= POS(2,4);
INST(17) <= INT_NUM(UNIDADES);
INST(18) <= BUCLE_FIN(1);

--INST() <= CODIGO_FIN(1);

-----------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------


end Behavioral;