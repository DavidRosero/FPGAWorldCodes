LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MotorPaP_Bipolar IS
		PORT( L_R, FS_HS: IN STD_LOGIC;
				CLK, RST, SPEED : IN STD_LOGIC;
				A, B, C, D: OUT STD_LOGIC;
				LED: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
				);
END MotorPaP_Bipolar;

--DECLARACIÓN DE VARIABLES
	
ARCHITECTURE BEHAVIORAL OF MotorPaP_Bipolar IS 
TYPE TYPE_STATE IS (S0,S1,S2,S3,S4,S5,S6,S7);
SIGNAL STATE: TYPE_STATE;
--DECLARACIÓN DE ESTADOS
SIGNAL AUX1, CLK1, AUX2, CLK2, VEL: STD_LOGIC;
SIGNAL COUNT1, COUNT2 :INTEGER:=1;
SIGNAL SALIDA : STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL X: STD_LOGIC_VECTOR (1 DOWNTO 0);

--DECLARACIÓN DE SEÑALES

BEGIN

VELOCIDAD_1HZ: PROCESS (CLK)
BEGIN
IF (CLK'EVENT AND CLK='1') THEN
		COUNT1 <= COUNT1+1;
		IF (COUNT1=25000000) THEN
			AUX1 <= NOT AUX1;
			COUNT1 <= 1;
		END IF;
	END IF;
END PROCESS;

CLK1 <= AUX1;
--DIVISOR DE FRECUENCIA A 1 HZ 

VELOCIDAD_500HZ: PROCESS (CLK)
BEGIN
	IF(CLK'EVENT AND CLK='1') THEN
			COUNT2 <= COUNT2+1;
			IF (COUNT2 = 50000) THEN
				AUX2 <= NOT AUX2;
				COUNT2 <= 1;
			END IF;
	END IF;
END PROCESS;
CLK2 <= AUX2;

--DIVISOR DE FRECUENCIA A 500 HZ

SEL_SPEED: PROCESS(CLK1,CLK2)
BEGIN
	IF (SPEED = '0') THEN	
		VEL <= CLK1;
		ELSE
			VEL <= CLK2;
			END IF;
		END PROCESS;
--SELECCCION DE LA VELOCIDAD DEL MOTOR
PROCESO_ESTADOS: PROCESS (RST, VEL)
BEGIN
X <= L_R&FS_HS;

--CONCATENACION DE LAS ENTRADAS L_R Y FS_HS (SENTIDO DE GIRO Y TIPO DE PASOS)

IF RST = '1' THEN
	STATE <= S0;
	--DECLARACIÓN DE ESTAD0 INICIAL
	
	ELSIF RISING_EDGE (VEL) THEN
	
CASE STATE IS 
	WHEN S0 =>
		IF (X = "00") THEN
		STATE <= S1;
		ELSIF (X = "01") THEN
		STATE <= S2;
		ELSIF (X = "10") THEN
		STATE <= S7;
		ELSIF (X = "11") THEN
		STATE <= S6;
		END IF;
	WHEN S1 =>
		IF (X = "00") THEN
		STATE <= S2;
		ELSIF (X = "01") THEN
		STATE <= S3;
		ELSIF (X = "10") THEN
		STATE <= S0;
		ELSIF (X = "11") THEN
		STATE <= S7;
		END IF;
	WHEN S2 =>
		IF (X = "00") THEN
		STATE <= S3;
		ELSIF (X = "01") THEN
		STATE <= S4;
		ELSIF (X = "10") THEN
		STATE <= S1;
		ELSIF (X = "11") THEN
		STATE <= S0;
		END IF;
	WHEN S3 =>
		IF (X = "00") THEN
		STATE <= S4;
		ELSIF (X = "01") THEN
		STATE <= S5;
		ELSIF (X = "10") THEN
		STATE <= S2;
		ELSIF (X = "11") THEN
		STATE <= S1;
		END IF;
	WHEN S4 =>
		IF (X = "00") THEN
		STATE <= S5;
		ELSIF (X = "01") THEN
		STATE <= S6;
		ELSIF (X = "10") THEN
		STATE <= S3;
		ELSIF (X = "11") THEN
		STATE <= S2;
		END IF;
	WHEN S5 =>
		IF (X = "00") THEN
		STATE <= S6;
		ELSIF (X = "01") THEN
		STATE <= S7;
		ELSIF (X = "10") THEN
		STATE <= S4;
		ELSIF (X = "11") THEN
		STATE <= S3;
		END IF;
	WHEN S6 =>
		IF (X = "00") THEN
		STATE <= S7;
		ELSIF (X = "01") THEN
		STATE <= S0;
		ELSIF (X = "10") THEN
		STATE <= S5;
		ELSIF (X = "11") THEN
		STATE <= S4;
		END IF;
	WHEN S7 =>
		IF (X = "00") THEN
		STATE <= S0;
		ELSIF (X = "01") THEN
		STATE <= S1;
		ELSIF (X = "10") THEN
		STATE <= S6;
		ELSIF (X = "11") THEN
		STATE <= S5;
		END IF;
	END CASE;
END IF;
END PROCESS;
--DEFINICIÓN DE CADA ESTADO CON SUS RESPECTIVAS CONDICIONES
LOGICA_SALIDA: PROCESS(STATE)
BEGIN

CASE STATE IS
	WHEN S0 => SALIDA <="0001";
	WHEN S1 => SALIDA <="0101";
	WHEN S2 => SALIDA <="0010";
	WHEN S3 => SALIDA <="1001";
	WHEN S4 => SALIDA <="1000";
	WHEN S5 => SALIDA <="1010";
	WHEN S6 => SALIDA <="0100";
	WHEN S7 => SALIDA <="0110";
END CASE;
END PROCESS;
--BLOQUE DE LA LOGICA DE SALIDA
SALIDAS_LEDS: PROCESS (CLK)
BEGIN
LED(0) <= SALIDA(0); 
LED(1) <= SALIDA(1);
LED(2) <= SALIDA(2);
LED(3) <= SALIDA(3);
END PROCESS;

A <= SALIDA(0); 
B <= SALIDA(1);
C <= SALIDA(2);
D <= SALIDA(3);

--ASIGNACION DE LAS VARIABLES DE SALIDA

END BEHAVIORAL;